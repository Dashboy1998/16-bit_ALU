package gate_delay is
	constant propagation: time := 10ns;
end gate_delay;